module  where


